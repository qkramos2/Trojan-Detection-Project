`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date: 10/05/2023 12:44:45 AM
// Design Name: 
// Module Name: wrapper
// Project Name: 
// Target Devices: 
// Tool Versions: 
// Description: 
// 
// Dependencies: 
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
//////////////////////////////////////////////////////////////////////////////////


module wrapper(
        in_val, 
        out_val
    );
    
input [177:0] in_val; 
output [122:0] out_val;


Circuit5315 wrap(

in_val[177],

in_val[176],

in_val[175],

in_val[174],

in_val[173],

in_val[172],

in_val[171],

in_val[170],

in_val[169],

in_val[168],

in_val[167],

in_val[166],

in_val[165],

in_val[164],

in_val[163],

in_val[162],

in_val[161],

in_val[160],

in_val[159],

in_val[158],

in_val[157],

in_val[156],

in_val[155],

in_val[154],

in_val[153],

in_val[152],

in_val[151],

in_val[150],

in_val[149],

in_val[148],

in_val[147],

in_val[146],

in_val[145],

in_val[144],

in_val[143],

in_val[142],

in_val[141],

in_val[140],

in_val[139],

in_val[138],

in_val[137],

in_val[136],

in_val[135],

in_val[134],

in_val[133],

in_val[132],

in_val[131],

in_val[130],

in_val[129],

in_val[128],

in_val[127],

in_val[126],

in_val[125],

in_val[124],

in_val[123],

in_val[122],

in_val[121],

in_val[120],

in_val[119],

in_val[118],

in_val[117],

in_val[116],

in_val[115],

in_val[114],

in_val[113],

in_val[112],

in_val[111],

in_val[110],

in_val[109],

in_val[108],

in_val[107],

in_val[106],

in_val[105],

in_val[104],

in_val[103],

in_val[102],

in_val[101],
in_val[100],

in_val[99],

in_val[98],

in_val[97],

in_val[96],

in_val[95],

in_val[94],

in_val[93],

in_val[92],

in_val[91],

in_val[90],

in_val[89],

in_val[88],

in_val[87],

in_val[86],

in_val[85],

in_val[84],

in_val[83],

in_val[82],

in_val[81],

in_val[80],

in_val[79],

in_val[78],

in_val[77],

in_val[76],

in_val[75],

in_val[74],

in_val[73],

in_val[72],

in_val[71],

in_val[70],

in_val[69],

in_val[68],

in_val[67],

in_val[66],

in_val[65],

in_val[64],

in_val[63],

in_val[62],

in_val[61],

in_val[60],

in_val[59],

in_val[58],

in_val[57],

in_val[56],

in_val[55],

in_val[54],

in_val[53],

in_val[52],

in_val[51],

in_val[50],

in_val[49],

in_val[48],

in_val[47],

in_val[46],

in_val[45],

in_val[44],

in_val[43],

in_val[42],

in_val[41],

in_val[40],
in_val[39],

in_val[38],

in_val[37],

in_val[36],

in_val[35],

in_val[34],

in_val[33],

in_val[32],

in_val[31],

in_val[30],

in_val[29],

in_val[28],

in_val[27],

in_val[26],

in_val[25],

in_val[24],

in_val[23],

in_val[22],

in_val[21],

in_val[20],

in_val[19],

in_val[18],

in_val[17],

in_val[16],

in_val[15],

in_val[14],

in_val[13],

in_val[12],

in_val[11],

in_val[10],

in_val[9],

in_val[8],

in_val[7],

in_val[6],

in_val[5],

in_val[4],

in_val[3],
in_val[2],

in_val[1],

in_val[0],
out_val[122],

out_val[121],

out_val[120],

out_val[119],

out_val[118],

out_val[117],

out_val[116],

out_val[115],

out_val[114],
out_val[113],

out_val[112],

out_val[111],

out_val[110],

out_val[109],

out_val[108],

out_val[107],

out_val[106],

out_val[105],

out_val[104],

out_val[103],

out_val[102],

out_val[101],

out_val[100],

out_val[99],

out_val[98],

out_val[97],

out_val[96],

out_val[95],

out_val[94],

out_val[93],

out_val[92],

out_val[91],

out_val[90],

out_val[89],

out_val[88],

out_val[87],

out_val[86],

out_val[85],

out_val[84],

out_val[83],

out_val[82],

out_val[81],

out_val[80],

out_val[79],

out_val[78],

out_val[77],

out_val[76],

out_val[75],

out_val[74],

out_val[73],

out_val[72],

out_val[71],

out_val[70],

out_val[69],

out_val[68],

out_val[67],

out_val[66],

out_val[65],

out_val[64],

out_val[63],

out_val[62],

out_val[61],

out_val[60],

out_val[59],

out_val[58],

out_val[57],

out_val[56],

out_val[55],

out_val[54],

out_val[53],

out_val[52],

out_val[51],

out_val[50],

out_val[49],

out_val[48],

out_val[47],

out_val[46],

out_val[45],

out_val[44],

out_val[43],

out_val[42],

out_val[41],

out_val[40],

out_val[39],

out_val[38],

out_val[37],

out_val[36],

out_val[35],

out_val[34],

out_val[33],

out_val[32],
out_val[31],

out_val[30],

out_val[29],

out_val[28],

out_val[27],

out_val[26],

out_val[25],

out_val[24],

out_val[23],

out_val[22],
out_val[21],

out_val[20],

out_val[19],

out_val[18],

out_val[17],

out_val[16],

out_val[15],

out_val[14],

out_val[13],

out_val[12],

out_val[11],

out_val[10],

out_val[9],

out_val[8],

out_val[7],

out_val[6],

out_val[5],

out_val[4],

out_val[3],

out_val[2],

out_val[1],

out_val[0]
);



endmodule
